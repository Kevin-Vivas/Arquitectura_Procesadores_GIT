module decodificador_hex(
  input wire A0,B0,C0,D0,
  output reg Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0
);

  always @(*) begin
    case({A0,B0,C0,D0})
      4'b0000: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b1000000; // 0
      4'b0001: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b1111001; // 1
      4'b0010: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0100100; // 2
      4'b0011: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0110000; // 3
      4'b0100: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0011001; // 4
      4'b0101: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0010010; // 5
      4'b0110: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0000010; // 6
      4'b0111: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b1111000; // 7
      4'b1000: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0000000; // 8
      4'b1001: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0010000; // 9
      4'b1010: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0001000; // A
      4'b1011: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0000011; // B
      4'b1100: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b1000110; // C
      4'b1101: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0100001; // D
      4'b1110: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0000110; // E
      4'b1111: {Aout0,Bout0,Cout0,Dout0,Eout0,Fout0,Gout0} = 7'b0001110; // F
    endcase
end

endmodule
